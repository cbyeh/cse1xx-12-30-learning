`timescale 1ns / 1ps

module my_and_gate(A,B,OUT);

	input A;
	input B;
	output OUT;
	
assign OUT = A&B;


endmodule