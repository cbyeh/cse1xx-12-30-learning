0 0 0 0 0 D11 D10 D9 <==  D8 D7 D6 D5 ...       D1

					   (D8) D7 D6 D5 ... D1 0									   10
																				   10
0 0 0 0 D11 D10 D9 D8					
					
																				  100
D11 D10 D09 D08 D07 D06 D05	 0
							 P8



							   <<
							   SC_out / SC_in